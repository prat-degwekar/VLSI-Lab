module bus(
	input [3:0]in,
	output out,
	input clk
);

assign out = in[0];
assign out = in[1];
assign out = in[2];
assign out = in[3];



endmodule
